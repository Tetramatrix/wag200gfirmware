time_zone=GMT+1 2 time_daylight= restore_default=0 wan_ifname=nas0 wan_mode=pppoe wan_iptype=Dynamic wan_ipaddr= wan_netmask= wan_gateway= wan_mtu=1500 wan_fix_dns=0 wan_dns1= wan_dns2= wan_macaddr= wan_encap=0 pppoa_encap=1 wan_vpivci_detect=1 wan_vpi=8 wan_vci=35 wan_account= wan_domain= wan_dod=1 wan_qos=ubr wan_pcr= wan_scr= wan_cmtu=auto dsl_modulation=MMODE dhcp_dns0= dhcp_dns1= dhcp_dns2= dhcp_wins= lan_if=br0 lan_ipaddr=192.168.1.1 lan_netmask=255.255.255.0 lan_bipaddr=192.168.1.255 dhcp_server_enable=1 dhcp_server_ip= dhcp_start_ip=192.168.1.100 dhcp_end_ip=192.168.1.149 dhcp_reserved= dhcp_lease=0 http_username=admin http_password=admin http_timeout=5 rt_static_route= rt_rip_version=1 rt_rip_direction=0 rt_rip_recvflag=1 rt_rip_sendflag=1 ddns_enable=0 ddns_service_provider=dyndns ddns_user_name= ddns_password= ddns_host_name= tzo_user_name= tzo_password= tzo_host_name= ddns_use_wildcards=0 pppoe_username= pppoe_password= pppoe_idle=5 pppoe_service= pppoe_redial=30 pppoa_username= pppoa_password= pppoa_ipaddr= wifi_ssid=linksys wifi_region= wifi_channel=11 wifi_auth_type=3 wifi_psk_pwd= wifi_psk_lifetime=3600 wifi_key_len=0 wifi_def_key=1 wifi_key1= wifi_key2= wifi_key3= wifi_key4= wifi_access_control=0 wifi_access_type=1 wifi_access_list= wifi_if_on=1 wifi_broadcast_ssid=1 wifi_wep_on=0 wifi_dot11_mode=0 wifi_dot11_iso=0 wifi_rate=0 wifi_radius_port=1812 wifi_beacon_period=100 wifi_dtim_period=1 wifi_rts=2347 wifi_frag=2346 mail_enable=0 mail_logfull=0 mail_sendlog=2 mail_server= mail_recipient= mail_dos=1 mail_portscan=1 mail_block=1 mail_sh_day=0 mail_sh_hour=1 log_dos=1 log_block=1 log_login=1 log_gateway=1 log_type=0 log_remote_ip= fw_nat=1 fw_block=1 fw_access_policy= fw_block_service=dns:17:53-53ping:1:0-0http:6:80-80https:6:443-443ftp:6:21-21pop3:6:110-110imap:6:143-143smtp:6:25-25nntp:6:119-119telnet:6:23-23snmp:17:161-161tftp:17:69-69ike:17:500-500 fw_block_trust_enable=0 fw_block_trust= fw_services_def=Any(ALL):any:1-65535Any(TCP):tcp:1-65535Any(UDP):udp:1-65535AIM:tcp:5190-5190BGP:tcp:179-179BOOTP_CLIENT:udp:68-68BOOTP_SERVER:udp:67-67CU-SEEME:both:7648-24032DNS:both:53-53FINGER:tcp:79-79FTP:tcp:20-21H.323:tcp:1720-1720HTTP:tcp:80-80HTTPS:tcp:443-443IDENT:tcp:113-113IRC:both:6667-6667NEWS:tcp:144-144NFS:udp:2049-2049NNTP:tcp:119-119RCMD:tcp:512-512REAL-AUDIO:tcp:7070-7070REXEC:tcp:514-514RLOGIN:tcp:513-513RTELNET:tcp:107-107RTSP:both:554-554SFTP:tcp:115-115SMTP:tcp:25-25SNMP:both:161-161SNMP-TRAPS:both:162-162SQL-NET:tcp:1521-1521SSH:both:22-22STRMWORKS:udp:1558-1558TACACS:udp:49-49TELNET:tcp:23-23TFTP:udp:69-69VDOLIVE:tcp:7000-7000VPN-IPSEC:udp:500-500VPN-L2TP:udp:1701-1701VPN-PPTP:tcp:1723-1723 fw_services= fw_in_rules=s:1:0:HTTP:0:0:80:80s:2:0:FTP:0:0:21:21s:3:0:FTP-Data:0:0:20:20s:4:0:Telnet:0:0:23:23s:5:0:SMTP:0:0:25:25s:6:0:TFTP:0:1:69:69s:7:0:finger:0:0:79:79s:8:0:NTP:0:1:123:123s:9:0:POP3:0:0:110:110s:10:0:NNTP:0:0:119:119s:11:0:SNMP:0:1:161:161s:12:0:CVS:0:0:2401:2401s:13:0:SMS:0:0:2701:2701s:14:0:SMS-rmctl:0:0:2702:2702 fw_out_rules= fw_dmz_enable=0 fw_dmz= fw_spi=1 fw_response_ping=0 fw_schedule=1111111:00:00-24:00 fw_time_zone=GMTb fw_remote=0 fw_remote_type= fw_remote_range_start= fw_remote_range_end= fw_remote_single= fw_remote_port=8080 ntp_custom=0 ntp_server= upnp_enable=1 upnp_adv_time=30 upnp_ttl=4 snmp_enable=0 snmp_read_community= snmp_set_community= snmp_sys_name= snmp_sys_contact= snmp_sys_location= snmp_trap_to= dhcpc_enable=1 ipsec_passthrough_enable=1 pppoe_passthrough_enable=1 pptp_passthrough_enable=1 l2tp_passthrough_enable=1 ping_size=60 ping_number=1 ping_interval=1000 ping_timeout=5000 fw_protection=1 fw_filter_proxy=0 fw_filter_cookies=0 fw_filter_java=0 fw_filter_activex=0 fw_block_wanrequest=1 log_enable=0 email_alert=0 dos_thresholds=20 smtp_mail_server= email_alert_addr= email_return_addr= qos_ds=disable qos_dslist=FTP:HHTTP:HTELNET:HSMTP:HPOP3:H0:L0:L0:L device_name=WAG200G lan_ifnames=br0 wlan0 language= igmp_proxy=1 wlan_mgr_enable=1 ipppoe_enable=0 timer_interval=3600  